module extender (
    input imm16, imm26,
    input extOp,
    output imm32
);
    
endmodule